n: 0 y:297889
n: 1 y:299526
n: 2 y:299094
