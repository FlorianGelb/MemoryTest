n: 0 y:298346
n: 1 y:299862
n: 2 y:296597
n: 0 y:299363
n: 0 y:299199
n: 0 y:297889
n: 1 y:299526
n: 2 y:299094
