n: 0 y:304040
n: 1 y:308040
n: 2 y:312040
n: 3 y:316040
n: 4 y:320040
n: 5 y:324040
n: 6 y:328040
n: 7 y:323904
n: 8 y:336040
n: 9 y:340040
n: 0 y:304040
n: 1 y:308040
n: 2 y:312040
n: 3 y:316040
n: 4 y:320040
n: 5 y:324040
n: 6 y:328040
n: 7 y:332040
n: 8 y:336040
n: 9 y:340040
n: 0 y:304040
n: 1 y:308040
n: 2 y:312040
n: 3 y:316040
n: 4 y:319448
n: 5 y:324040
n: 6 y:324456
n: 0 y:304040
n: 1 y:308040
n: 2 y:312040
n: 3 y:316040
n: 4 y:311904
n: 5 y:324040
n: 6 y:328040
n: 7 y:332040
n: 8 y:334024
n: 9 y:331904
n: 0 y:300240
n: 1 y:308040
n: 2 y:312040
n: 3 y:309512
n: 4 y:314808
n: 5 y:322640
n: 6 y:325952
n: 7 y:330640
n: 8 y:335688
n: 9 y:338528
n: 10 y:344056
n: 11 y:339920
n: 12 y:352016
n: 13 y:353760
n: 14 y:354824
n: 15 y:363328
n: 16 y:359920
n: 17 y:363920
n: 18 y:369624
n: 19 y:371920
n: 20 y:382656
n: 21 y:379920
n: 22 y:389856
n: 23 y:393760
n: 24 y:398736
n: 25 y:395920
n: 26 y:408016
n: 27 y:412056
n: 28 y:416056
n: 29 y:416256
n: 30 y:415920
n: 31 y:419920
n: 32 y:432056
n: 33 y:436056
n: 34 y:440056
n: 35 y:444056
n: 36 y:448056
n: 37 y:448424
n: 38 y:454448
n: 39 y:452016
n: 40 y:464056
n: 41 y:468056
n: 42 y:472056
n: 43 y:467920
n: 44 y:480056
n: 45 y:484056
n: 46 y:488056
n: 47 y:491696
n: 48 y:496016
n: 49 y:500056
n: 50 y:504056
n: 51 y:507424
n: 52 y:503920
n: 53 y:515424
n: 54 y:520056
n: 55 y:515920
n: 56 y:528056
n: 57 y:532056
n: 58 y:536056
n: 59 y:531920
n: 60 y:544056
n: 61 y:548056
n: 62 y:1225512
n: 63 y:547920
n: 64 y:551920
n: 65 y:555920
n: 66 y:568056
n: 67 y:570712
n: 68 y:567976
n: 69 y:579384
n: 70 y:584112
n: 71 y:579976
n: 72 y:587984
n: 73 y:594752
n: 74 y:598504
n: 75 y:595976
n: 76 y:599976
n: 77 y:603976
n: 78 y:607976
n: 79 y:620112
n: 80 y:624112
n: 81 y:628112
n: 82 y:623976
n: 83 y:636112
n: 84 y:640112
n: 85 y:644112
n: 86 y:648112
n: 87 y:647624
n: 88 y:656072
n: 89 y:651976
n: 90 y:655976
n: 91 y:668112
n: 92 y:672072
n: 93 y:667976
n: 94 y:680112
n: 95 y:675976
n: 96 y:688112
n: 97 y:691800
n: 98 y:687976
n: 99 y:691976
n: 100 y:695976
n: 101 y:708112
n: 102 y:703976
n: 103 y:716112
n: 104 y:711976
n: 105 y:718784
n: 106 y:719976
n: 107 y:723976
n: 108 y:727976
n: 109 y:731976
n: 110 y:744112
n: 111 y:747480
n: 112 y:752112
n: 113 y:756112
n: 114 y:760112
n: 115 y:296864
n: 116 y:768112
n: 117 y:771520
n: 118 y:776112
n: 119 y:303768
n: 120 y:784112
n: 121 y:296040
n: 122 y:783976
n: 123 y:295944
n: 124 y:304080
n: 125 y:804112
n: 126 y:799976
n: 127 y:298920
n: 128 y:304080
n: 129 y:303768
n: 130 y:304080
n: 131 y:302720
n: 132 y:295944
n: 133 y:295944
n: 134 y:295944
n: 135 y:303768
n: 136 y:295944
n: 137 y:299728
n: 138 y:295944
n: 139 y:295944
n: 140 y:299704
n: 141 y:300008
n: 142 y:295944
n: 143 y:304080
n: 144 y:298960
n: 145 y:300704
n: 146 y:295944
n: 147 y:300008
n: 148 y:295944
n: 149 y:295944
n: 150 y:303768
n: 151 y:301376
n: 152 y:302608
n: 153 y:295944
n: 154 y:302720
n: 155 y:304080
n: 156 y:302720
n: 157 y:304080
n: 158 y:304080
n: 159 y:304080
n: 160 y:304080
n: 161 y:303448
n: 162 y:295944
n: 163 y:303448
n: 164 y:304080
n: 165 y:295944
n: 166 y:303488
n: 167 y:295944
n: 168 y:295944
n: 169 y:304080
n: 170 y:295944
n: 171 y:295944
n: 172 y:295944
n: 173 y:295944
n: 174 y:295944
n: 175 y:304080
n: 176 y:302720
n: 177 y:301880
n: 178 y:304080
n: 179 y:300320
n: 180 y:304080
n: 181 y:303448
n: 182 y:295944
n: 183 y:295944
n: 184 y:300320
n: 185 y:303488
n: 186 y:303448
n: 187 y:295944
n: 188 y:297552
n: 189 y:295944
n: 190 y:303448
n: 191 y:295944
n: 192 y:304080
n: 193 y:295944
n: 194 y:296864
n: 195 y:296864
n: 196 y:303768
n: 197 y:295944
n: 198 y:304080
n: 199 y:296864
n: 200 y:295944
n: 201 y:295944
n: 202 y:295944
n: 203 y:295944
n: 204 y:303768
n: 205 y:300008
n: 206 y:303488
n: 207 y:295944
n: 208 y:299664
n: 209 y:295944
n: 210 y:303768
n: 211 y:295944
n: 212 y:304080
n: 213 y:295944
n: 214 y:298752
n: 215 y:303488
n: 216 y:302512
n: 217 y:295944
n: 218 y:300488
n: 219 y:295944
n: 220 y:300008
n: 221 y:303488
n: 222 y:304080
n: 223 y:304080
n: 224 y:303448
n: 225 y:295944
n: 226 y:301784
n: 227 y:295944
n: 228 y:295944
n: 229 y:303488
n: 230 y:304080
n: 231 y:295944
n: 232 y:298752
n: 233 y:295944
n: 234 y:304080
n: 235 y:295944
n: 236 y:298752
n: 237 y:302680
n: 238 y:300320
n: 239 y:295944
n: 240 y:297552
n: 241 y:295944
n: 242 y:302720
n: 243 y:303768
n: 244 y:303768
n: 245 y:304080
n: 246 y:295944
n: 247 y:295944
n: 248 y:302512
n: 249 y:295944
n: 250 y:298864
n: 251 y:295944
n: 252 y:295944
n: 253 y:303768
n: 254 y:302512
n: 255 y:304080
n: 256 y:295944
n: 257 y:295944
n: 258 y:295944
n: 259 y:304080
n: 260 y:302680
n: 261 y:295944
n: 262 y:295944
n: 263 y:295944
n: 264 y:295944
n: 265 y:298472
n: 266 y:304080
n: 267 y:300648
n: 268 y:301728
n: 269 y:302512
n: 270 y:295944
n: 271 y:304080
n: 272 y:303768
n: 273 y:295944
n: 274 y:304080
n: 275 y:295944
n: 276 y:304080
n: 277 y:295944
n: 278 y:295944
n: 279 y:303488
n: 280 y:303768
n: 281 y:303768
n: 282 y:295944
n: 283 y:298376
n: 284 y:304080
n: 285 y:303768
n: 286 y:304080
n: 287 y:295944
n: 288 y:295944
n: 289 y:295944
n: 290 y:295944
n: 291 y:304080
n: 292 y:295944
n: 293 y:303768
n: 294 y:295944
n: 295 y:303768
n: 296 y:302720
n: 297 y:299704
n: 298 y:295944
n: 299 y:298472
n: 300 y:299824
n: 301 y:295944
n: 302 y:304080
n: 303 y:300416
n: 304 y:298960
n: 305 y:304080
n: 306 y:295944
n: 307 y:295944
n: 308 y:303768
n: 309 y:298752
n: 310 y:304080
n: 311 y:302720
n: 312 y:304080
n: 313 y:295944
n: 314 y:295944
n: 315 y:295944
n: 316 y:304080
n: 317 y:303768
n: 318 y:300320
n: 319 y:304080
n: 320 y:303768
n: 321 y:295944
n: 322 y:303488
n: 323 y:295944
n: 324 y:295944
n: 325 y:295944
n: 326 y:302512
n: 327 y:303488
n: 328 y:300008
n: 329 y:298752
n: 330 y:297688
n: 331 y:296960
n: 332 y:299728
n: 333 y:295944
n: 334 y:298752
n: 335 y:302064
n: 336 y:1648096
n: 337 y:303768
n: 338 y:304080
n: 339 y:297688
n: 340 y:304080
n: 341 y:304080
n: 342 y:295944
n: 343 y:295944
n: 344 y:303768
n: 345 y:304080
n: 346 y:295944
n: 347 y:295944
n: 348 y:295944
n: 349 y:304080
n: 350 y:304080
n: 351 y:295944
n: 352 y:295944
n: 353 y:297552
n: 354 y:295944
n: 355 y:295944
n: 356 y:302064
n: 357 y:295944
n: 358 y:295944
n: 359 y:303488
n: 360 y:295944
n: 361 y:304080
n: 362 y:295944
n: 363 y:303448
n: 364 y:302720
n: 365 y:295944
n: 366 y:295944
n: 367 y:303448
n: 368 y:295944
n: 369 y:303768
n: 370 y:304080
n: 371 y:302680
n: 372 y:295944
n: 373 y:295944
n: 374 y:304080
n: 375 y:303448
n: 376 y:295944
n: 377 y:304080
n: 378 y:304080
n: 379 y:303768
n: 380 y:295944
n: 381 y:295944
n: 382 y:304080
n: 383 y:299728
n: 384 y:304080
n: 385 y:295944
n: 386 y:295944
n: 387 y:295944
n: 388 y:303488
n: 389 y:302608
n: 390 y:304080
n: 391 y:302720
n: 392 y:303768
n: 393 y:304080
n: 394 y:295944
n: 395 y:298752
n: 396 y:303768
n: 397 y:295944
n: 398 y:303488
n: 399 y:300768
n: 400 y:295944
n: 401 y:295944
n: 402 y:301472
n: 403 y:295944
n: 404 y:304080
n: 405 y:304080
n: 406 y:296864
n: 407 y:300320
n: 408 y:304080
n: 409 y:298848
n: 410 y:304080
n: 411 y:303768
n: 412 y:298432
n: 413 y:304080
n: 414 y:295944
n: 415 y:295944
n: 416 y:301240
n: 417 y:303768
n: 418 y:295944
n: 419 y:295944
n: 420 y:304080
n: 421 y:295944
n: 422 y:303448
n: 423 y:295944
n: 424 y:304080
n: 425 y:304080
n: 426 y:303768
n: 427 y:295944
n: 428 y:295944
n: 429 y:295944
n: 430 y:298960
n: 431 y:295944
n: 432 y:295944
n: 433 y:299824
n: 434 y:303448
n: 435 y:295944
n: 436 y:303768
n: 437 y:295944
n: 438 y:295944
n: 439 y:304080
n: 440 y:299592
n: 441 y:298960
n: 442 y:304080
n: 443 y:303448
n: 444 y:295944
n: 445 y:295944
n: 446 y:295944
n: 447 y:295944
n: 448 y:304080
n: 449 y:295944
n: 450 y:298848
n: 451 y:304080
n: 452 y:295944
n: 453 y:301144
n: 454 y:301880
n: 455 y:304080
n: 456 y:300008
n: 457 y:303488
n: 458 y:302608
n: 459 y:297688
n: 460 y:295944
n: 461 y:304080
n: 462 y:304080
n: 463 y:304080
n: 464 y:302512
n: 465 y:303352
n: 466 y:295944
n: 467 y:304080
n: 468 y:303768
n: 469 y:303488
n: 470 y:304080
n: 471 y:304080
n: 472 y:295944
n: 473 y:304080
n: 474 y:295944
n: 475 y:2196056
n: 476 y:295944
n: 477 y:300704
n: 478 y:300008
n: 479 y:304080
n: 480 y:303488
n: 481 y:298960
n: 482 y:295944
n: 483 y:295944
n: 484 y:295944
n: 485 y:303488
n: 486 y:302608
n: 487 y:302608
n: 488 y:297688
n: 489 y:303768
n: 490 y:304080
n: 491 y:304080
n: 492 y:297688
n: 493 y:302512
n: 494 y:295944
n: 495 y:296728
n: 496 y:300488
n: 497 y:295944
n: 498 y:304080
n: 499 y:295944
n: 500 y:302720
n: 501 y:295944
n: 502 y:304080
n: 503 y:303448
n: 504 y:304080
n: 505 y:295944
n: 506 y:295944
n: 507 y:304080
n: 508 y:304080
n: 509 y:304080
n: 510 y:303728
n: 511 y:304080
n: 512 y:304080
n: 513 y:295944
n: 514 y:298752
n: 515 y:2364096
n: 516 y:297648
n: 517 y:2363960
n: 518 y:2367960
n: 519 y:295944
n: 520 y:303768
n: 521 y:2385800
n: 522 y:295944
n: 523 y:295944
n: 524 y:304080
n: 525 y:2402080
n: 526 y:304080
n: 527 y:304080
n: 528 y:298848
n: 529 y:304080
n: 530 y:302512
n: 531 y:2428096
n: 532 y:304080
n: 533 y:297592
n: 534 y:298960
n: 535 y:297744
n: 536 y:295944
n: 537 y:298960
n: 538 y:2456096
n: 539 y:300320
n: 540 y:2455960
n: 541 y:2459960
n: 542 y:2470488
n: 543 y:2476096
n: 544 y:304080
n: 545 y:298960
n: 546 y:296768
n: 547 y:304080
n: 548 y:304080
n: 549 y:303488
n: 550 y:299704
n: 551 y:304080
n: 552 y:2511464
n: 553 y:304080
n: 554 y:2511960
n: 555 y:2524096
n: 556 y:2527784
n: 557 y:304080
n: 558 y:2535744
n: 559 y:299704
n: 560 y:304080
n: 561 y:2546776
n: 562 y:303768
n: 563 y:2556096
n: 564 y:295944
n: 565 y:2560512
n: 566 y:2568096
n: 567 y:295944
n: 568 y:2576096
n: 569 y:295944
n: 570 y:2584096
n: 571 y:304080
n: 572 y:295944
n: 573 y:2587960
n: 574 y:2591960
n: 575 y:2604096
n: 576 y:2608096
n: 577 y:2603960
n: 578 y:2616096
n: 579 y:2619464
n: 580 y:300008
n: 581 y:302720
n: 582 y:2623960
n: 583 y:2636096
n: 584 y:2631960
n: 585 y:2635960
n: 586 y:303448
n: 587 y:2650008
n: 588 y:2655056
n: 589 y:304080
n: 590 y:2655960
n: 591 y:304080
n: 592 y:2672096
n: 593 y:2674528
n: 594 y:2671960
n: 595 y:302720
n: 596 y:2679960
n: 597 y:304080
n: 598 y:2688784
n: 599 y:2698080
n: 600 y:2695960
n: 601 y:304080
n: 602 y:2710528
n: 603 y:2707960
n: 604 y:2719056
n: 605 y:2723504
n: 606 y:2728096
n: 607 y:2732056
n: 608 y:2736096
n: 609 y:295944
n: 610 y:2743464
n: 611 y:2748096
n: 612 y:2747664
n: 613 y:2747960
n: 614 y:2759744
n: 615 y:2764096
n: 616 y:2764024
n: 617 y:2772096
n: 618 y:2776096
n: 619 y:2778080
n: 620 y:2775960
n: 621 y:2788096
n: 622 y:2790528
n: 623 y:2796096
n: 624 y:2791960
n: 625 y:2803784
n: 626 y:2808096
n: 627 y:2805608
n: 628 y:2813800
n: 629 y:304080
n: 630 y:2823504
n: 631 y:2827464
n: 632 y:2829800
n: 633 y:2834736
n: 634 y:2831960
n: 635 y:2844096
n: 636 y:2846528
n: 637 y:2852096
n: 638 y:2847960
n: 639 y:2851960
n: 640 y:2855960
n: 641 y:2859960
n: 642 y:304080
n: 643 y:2876096
n: 644 y:2880096
n: 645 y:2875960
n: 646 y:2887464
n: 647 y:2883960
n: 648 y:2887960
n: 649 y:2900096
n: 650 y:2903784
n: 651 y:2908096
n: 652 y:2910080
n: 653 y:2907960
n: 654 y:2917952
n: 655 y:2923784
n: 656 y:2922992
n: 657 y:2931784
n: 658 y:2928784
n: 659 y:295944
n: 660 y:2944096
n: 661 y:2948096
n: 662 y:2952096
n: 663 y:2947960
n: 664 y:298752
n: 665 y:2964096
n: 666 y:2968096
n: 667 y:2972096
n: 668 y:2976096
n: 669 y:2971960
n: 670 y:2984096
n: 671 y:2986696
n: 672 y:2986768
n: 673 y:2996096
n: 674 y:2997744
n: 675 y:3001896
n: 676 y:2999960
n: 677 y:3003960
n: 678 y:298752
n: 679 y:3011960
n: 680 y:295944
n: 681 y:3023744
n: 682 y:3023960
n: 683 y:3027960
n: 684 y:3039744
n: 685 y:3040664
n: 686 y:3048096
n: 687 y:3052096
n: 688 y:295944
n: 689 y:3051960
n: 690 y:3055960
n: 691 y:3059960
n: 692 y:3064976
n: 693 y:3076096
n: 694 y:295944
n: 695 y:3083784
n: 696 y:3079960
n: 697 y:3092096
n: 698 y:3087960
n: 699 y:295944
n: 700 y:3104096
n: 701 y:3108096
n: 702 y:3112096
n: 703 y:3116096
n: 704 y:3119464
n: 705 y:3122528
n: 706 y:3128096
n: 707 y:3126768
n: 708 y:3127960
n: 709 y:3137800
n: 710 y:3138976
n: 711 y:3142768
n: 712 y:3151464
n: 713 y:3147960
n: 714 y:3160096
n: 715 y:3164096
n: 716 y:3167504
n: 717 y:3170528
n: 718 y:3167960
n: 719 y:3174976
n: 720 y:3180464
n: 721 y:3188096
n: 722 y:3192096
n: 723 y:3187960
n: 724 y:3196432
n: 725 y:3195960
n: 726 y:3205160
n: 727 y:3212096
n: 728 y:3216096
n: 729 y:295944
n: 730 y:3224096
n: 731 y:3219960
n: 732 y:3232096
n: 733 y:3230864
n: 734 y:3231960
n: 735 y:3244096
n: 736 y:3239960
n: 737 y:3243960
n: 738 y:3247960
n: 739 y:3258488
n: 740 y:3262080
n: 741 y:3268096
n: 742 y:3263960
n: 743 y:3276096
n: 744 y:3280096
n: 745 y:3282488
n: 746 y:3286008
n: 747 y:3288512
n: 748 y:3287960
n: 749 y:3291960
n: 750 y:3302008
n: 751 y:3307464
n: 752 y:3306768
n: 753 y:295944
n: 754 y:3320096
n: 755 y:3315960
n: 756 y:3319960
n: 757 y:3323960
n: 758 y:3334488
n: 759 y:3331960
n: 760 y:3335960
n: 761 y:3339960
n: 762 y:3343960
n: 763 y:3347960
n: 764 y:3358008
n: 765 y:3355960
n: 766 y:3359960
n: 767 y:3372096
n: 768 y:3367960
n: 769 y:3378488
n: 770 y:3375960
n: 771 y:3387504
n: 772 y:3383960
n: 773 y:3394080
n: 774 y:3391960
n: 775 y:3395960
n: 776 y:3408096
n: 777 y:3403960
n: 778 y:3414008
n: 779 y:3420096
n: 780 y:3415960
n: 781 y:3428096
n: 782 y:3432096
n: 783 y:3436096
n: 784 y:3431960
n: 785 y:3444096
n: 786 y:3448096
n: 787 y:3448024
n: 788 y:3451704
n: 789 y:3451960
n: 790 y:3455960
n: 791 y:3468096
n: 792 y:3471784
n: 793 y:3475504
n: 794 y:3478736
n: 795 y:3475960
n: 796 y:3481608
n: 797 y:3483960
n: 798 y:3496096
n: 799 y:3500096
n: 800 y:3495960
n: 801 y:3507744
n: 802 y:3509896
n: 803 y:3514736
n: 804 y:3519784
n: 805 y:3518976
n: 806 y:3527784
n: 807 y:3532096
n: 808 y:3536096
n: 809 y:3540096
n: 810 y:3544056
n: 811 y:3548096
n: 812 y:3543960
n: 813 y:3556096
n: 814 y:3553608
n: 815 y:3563784
n: 816 y:3564432
n: 817 y:3570528
n: 818 y:3576096
n: 819 y:3571960
n: 820 y:3584096
n: 821 y:3588096
n: 822 y:3592096
n: 823 y:3587960
n: 824 y:3591960
n: 825 y:3595960
n: 826 y:3599960
n: 827 y:3612096
n: 828 y:3614528
n: 829 y:3616512
n: 830 y:3619984
n: 831 y:3619960
n: 832 y:3631744
n: 833 y:3630768
n: 834 y:3631960
n: 835 y:3641952
n: 836 y:3639960
n: 837 y:3644880
n: 838 y:3652336
n: 839 y:3654352
n: 840 y:3664096
n: 841 y:3665488
n: 842 y:3663960
n: 843 y:3671720
n: 844 y:3675984
n: 845 y:3683368
n: 846 y:3679960
n: 847 y:3688336
n: 848 y:3687960
n: 849 y:3697952
n: 850 y:3697472
n: 851 y:3706584
n: 852 y:3712096
n: 853 y:3716096
n: 854 y:3720096
n: 855 y:3715960
n: 856 y:3726008
n: 857 y:3732096
n: 858 y:3727960
n: 859 y:3731960
n: 860 y:3735960
n: 861 y:3748096
n: 862 y:3743960
n: 863 y:3755056
n: 864 y:3751960
n: 865 y:3762080
n: 866 y:3759960
n: 867 y:3763960
n: 868 y:3770768
n: 869 y:3780096
n: 870 y:3784096
n: 871 y:3779960
n: 872 y:3783960
n: 873 y:3796096
n: 874 y:3791960
n: 875 y:3802488
n: 876 y:3808096
n: 877 y:3812096
n: 878 y:3814528
n: 879 y:3820096
n: 880 y:3815960
n: 881 y:3819960
n: 882 y:3823960
n: 883 y:3831984
n: 884 y:3834768
n: 885 y:3844096
n: 886 y:3839960
n: 887 y:3852096
n: 888 y:3847960
n: 889 y:3858584
n: 890 y:3862696
n: 891 y:3867784
n: 892 y:3870736
n: 893 y:3876096
n: 894 y:3880096
n: 895 y:3883784
n: 896 y:3886736
n: 897 y:3883960
n: 898 y:3891664
n: 899 y:3900096
n: 900 y:3895960
n: 901 y:3908096
n: 902 y:3912096
n: 903 y:3913896
n: 904 y:3917744
n: 905 y:3915960
n: 906 y:3928096
n: 907 y:3924936
n: 908 y:3927960
n: 909 y:3931960
n: 910 y:3943464
n: 911 y:3948096
n: 912 y:3944880
n: 913 y:3954736
n: 914 y:3951960
n: 915 y:3958488
n: 916 y:3967784
n: 917 y:3967984
n: 918 y:3975784
n: 919 y:3978008
n: 920 y:3975960
n: 921 y:3979960
n: 922 y:3990488
n: 923 y:3987960
n: 924 y:4000096
n: 925 y:3996056
n: 926 y:4007464
n: 927 y:4010736
n: 928 y:4016096
n: 929 y:4011960
n: 930 y:4024096
n: 931 y:4019960
n: 932 y:4032096
n: 933 y:4027960
n: 934 y:4031960
n: 935 y:4042696
n: 936 y:4048096
n: 937 y:4052096
n: 938 y:4047960
n: 939 y:4060096
n: 940 y:4055960
n: 941 y:4068096
n: 942 y:4063960
n: 943 y:4076096
n: 944 y:4079784
n: 945 y:4080528
n: 946 y:4087464
n: 947 y:4092096
n: 948 y:4090992
n: 949 y:4093608
n: 950 y:4104096
n: 951 y:4108096
n: 952 y:4112096
n: 953 y:4107960
n: 954 y:4119784
n: 955 y:4115960
n: 956 y:4126080
n: 957 y:4132096
n: 958 y:4136096
n: 959 y:4140096
n: 960 y:4141984
n: 961 y:4139960
n: 962 y:4144976
n: 963 y:4154736
n: 964 y:4155800
n: 965 y:4155960
n: 966 y:4168096
n: 967 y:4163960
n: 968 y:4167960
n: 969 y:4178584
n: 970 y:4175960
n: 971 y:4179960
n: 972 y:4190488
n: 973 y:4196096
n: 974 y:4191960
n: 975 y:4204096
n: 976 y:4206736
n: 977 y:4209800
n: 978 y:4207960
n: 979 y:4211960
n: 980 y:4224096
n: 981 y:4223608
n: 982 y:4232096
n: 983 y:4234584
n: 984 y:4239784
n: 985 y:4235960
n: 986 y:4248096
n: 987 y:4243960
n: 988 y:4255368
n: 989 y:4258736
n: 990 y:4259608
n: 991 y:4259960
n: 992 y:4271744
n: 993 y:4275744
n: 994 y:4271960
n: 995 y:4275960
n: 996 y:4288096
n: 997 y:4291504
n: 998 y:4296096
n: 999 y:4300096
n: 0 y:296000
n: 1 y:308040
n: 2 y:312040
n: 3 y:316040
n: 4 y:320040
n: 5 y:324040
n: 6 y:328040
n: 7 y:332000
n: 8 y:336040
n: 9 y:340040
n: 0 y:300240
n: 1 y:308040
n: 2 y:311728
n: 3 y:316040
n: 4 y:320040
n: 5 y:324040
n: 6 y:328040
n: 7 y:326880
n: 8 y:336040
n: 9 y:340040
n: 0 y:302720
n: 1 y:303928
n: 2 y:311728
n: 3 y:316040
n: 4 y:320000
n: 5 y:324040
n: 6 y:328040
n: 7 y:332040
n: 8 y:336040
n: 9 y:339448
n: 10 y:335920
n: 11 y:347016
n: 12 y:352056
n: 13 y:356056
n: 14 y:360056
n: 15 y:364056
n: 16 y:368056
n: 17 y:372056
n: 18 y:376056
n: 19 y:380056
n: 20 y:380296
n: 21 y:388056
n: 22 y:391328
n: 23 y:396056
n: 24 y:400056
n: 25 y:404056
n: 26 y:408056
n: 27 y:409120
n: 28 y:416056
n: 29 y:420056
n: 30 y:424056
n: 31 y:428056
n: 32 y:432056
n: 33 y:436056
n: 34 y:440056
n: 35 y:444016
n: 36 y:448016
n: 37 y:452056
n: 38 y:456056
n: 39 y:451920
n: 40 y:464056
n: 41 y:468056
n: 42 y:472016
n: 43 y:475744
n: 44 y:471920
n: 45 y:483424
n: 46 y:486696
n: 47 y:492056
n: 48 y:489568
n: 49 y:495568
n: 0 y:296688
n: 1 y:304048
n: 2 y:304048
n: 3 y:302368
n: 4 y:303704
n: 5 y:295928
n: 6 y:302664
n: 7 y:295936
n: 8 y:301928
n: 9 y:295944
n: 10 y:300608
n: 11 y:298760
n: 12 y:303776
n: 13 y:304096
n: 14 y:303464
n: 15 y:304104
n: 16 y:304104
n: 17 y:304112
n: 18 y:295976
n: 19 y:295984
n: 20 y:304120
n: 21 y:304128
n: 22 y:295992
n: 23 y:304136
n: 24 y:303824
n: 25 y:303512
n: 26 y:304144
n: 27 y:304152
n: 28 y:304152
n: 29 y:304160
n: 30 y:304160
n: 31 y:304168
n: 32 y:304168
n: 33 y:304176
n: 34 y:296040
n: 35 y:304184
n: 36 y:296048
n: 37 y:296056
n: 38 y:296056
n: 39 y:304200
n: 40 y:296064
n: 41 y:296072
n: 42 y:302640
n: 43 y:296080
n: 44 y:298984
n: 45 y:304224
n: 46 y:302072
n: 47 y:302144
n: 48 y:296096
n: 49 y:296104
n: 0 y:304040
n: 1 y:304048
n: 2 y:303416
n: 0 y:303688
n: 1 y:304048
n: 2 y:295912
n: 3 y:295920
n: 4 y:302736
n: 5 y:302664
n: 6 y:299672
n: 7 y:300640
n: 8 y:302464
n: 9 y:298752
n: 10 y:303352
n: 11 y:302480
n: 12 y:304088
n: 13 y:302008
n: 14 y:303744
n: 15 y:295968
n: 16 y:295968
n: 17 y:302504
n: 18 y:300000
n: 19 y:301920
n: 20 y:300008
n: 21 y:302520
n: 22 y:301832
n: 23 y:302624
n: 24 y:303504
n: 25 y:301848
n: 26 y:302536
n: 27 y:298824
n: 28 y:296016
n: 29 y:302648
n: 30 y:302760
n: 31 y:302560
n: 32 y:296032
n: 33 y:299056
n: 34 y:299056
n: 35 y:297696
n: 36 y:296048
n: 37 y:302584
n: 38 y:298864
n: 39 y:296064
n: 40 y:304200
n: 41 y:304208
n: 42 y:303616
n: 43 y:304136
n: 44 y:304216
n: 45 y:304224
n: 46 y:304224
n: 47 y:304232
n: 48 y:304232
n: 49 y:304240
n: 0 y:301840
n: 1 y:303696
n: 2 y:295912
n: 3 y:301760
n: 4 y:304056
n: 5 y:304064
n: 6 y:300264
n: 7 y:298424
n: 8 y:304072
n: 9 y:295944
n: 10 y:295944
n: 11 y:295952
n: 12 y:295952
n: 13 y:304096
n: 14 y:304096
n: 15 y:304104
n: 16 y:295968
n: 17 y:295976
n: 18 y:302752
n: 19 y:303448
n: 20 y:300008
n: 21 y:295992
n: 22 y:303816
n: 23 y:296000
n: 24 y:304136
n: 25 y:302744
n: 26 y:299848
n: 27 y:296936
n: 28 y:302752
n: 29 y:304160
n: 30 y:303528
n: 31 y:298952
n: 32 y:303496
n: 33 y:302568
n: 34 y:303448
n: 35 y:302864
n: 36 y:296048
n: 37 y:301216
n: 38 y:302680
n: 39 y:304200
n: 40 y:302800
n: 41 y:296072
n: 42 y:300544
n: 43 y:304216
n: 44 y:296080
n: 45 y:298896
n: 46 y:296184
n: 47 y:296096
n: 48 y:299112
n: 49 y:299008
n: 0 y:295904
n: 1 y:302688
n: 2 y:303008
n: 3 y:303328
n: 4 y:303744
n: 5 y:304024
n: 6 y:304064
n: 7 y:296760
n: 8 y:303760
n: 9 y:302472
n: 10 y:304080
n: 11 y:304088
n: 12 y:304048
n: 13 y:302736
n: 14 y:301216
n: 15 y:303376
n: 16 y:304104
n: 17 y:304072
n: 18 y:304112
n: 19 y:304120
n: 20 y:299000
n: 21 y:304128
n: 22 y:304128
n: 23 y:304136
n: 24 y:304136
n: 25 y:304144
n: 26 y:303832
n: 27 y:304152
n: 28 y:300040
n: 29 y:296024
n: 30 y:297768
n: 31 y:296032
n: 32 y:303856
n: 33 y:304176
n: 34 y:304176
n: 35 y:302824
n: 36 y:302168
n: 37 y:304192
n: 38 y:304192
n: 39 y:304200
n: 40 y:303608
n: 41 y:303576
n: 42 y:304208
n: 43 y:304216
n: 44 y:303488
n: 45 y:304224
n: 46 y:304224
n: 47 y:296096
n: 48 y:304232
n: 49 y:304240
n: 0 y:303920.0
n: 1 y:299588.8
n: 2 y:300391.2
n: 3 y:300624.0
n: 4 y:300844.8
n: 5 y:302044.0
n: 6 y:302149.6
n: 7 y:300774.4
n: 8 y:303454.4
n: 9 y:302170.4
n: 10 y:303023.2
n: 11 y:301084.0
n: 12 y:303246.4
n: 13 y:300303.2
n: 14 y:303293.6
n: 15 y:303047.2
n: 16 y:303507.2
n: 17 y:302745.6
n: 18 y:302699.2
n: 19 y:302516.0
n: 20 y:303576.0
n: 21 y:302334.4
n: 22 y:303110.4
n: 23 y:302285.6
n: 24 y:303580.8
n: 25 y:301772.8
n: 26 y:301475.2
n: 27 y:300174.4
n: 28 y:302800.8
n: 29 y:303769.6
n: 30 y:301240.0
n: 31 y:302052.8
n: 32 y:300784.0
n: 33 y:302952.0
n: 34 y:302744.0
n: 35 y:304060.0
n: 36 y:304060.0
n: 37 y:304024.8
n: 38 y:303297.6
n: 39 y:301515.2
n: 40 y:301584.0
n: 41 y:302741.6
n: 42 y:303696.8
n: 43 y:301049.6
n: 44 y:301555.2
n: 45 y:299882.4
n: 46 y:303636.8
n: 47 y:303058.4
n: 48 y:303215.2
n: 49 y:303044.8
n: 0 y:297566
n: 1 y:298706
n: 2 y:301531
n: 0 y:303006
n: 1 y:303965
n: 2 y:302978
n: 0 y:302986
n: 1 y:302708
n: 2 y:302120
n: 0 y:297889
n: 1 y:299526
n: 2 y:299094
n: 0 y:296349
n: 1 y:339732
n: 2 y:379231
n: 3 y:419348
n: 4 y:458149
n: 5 y:498926
n: 6 y:540396
n: 7 y:549466
n: 8 y:617003
n: 9 y:657637
n: 10 y:618124
n: 11 y:651103
n: 12 y:634204
n: 13 y:348739
n: 14 y:352511
n: 15 y:296224
n: 16 y:295944
n: 17 y:296032
n: 18 y:296224
n: 19 y:372120
n: 20 y:295944
n: 21 y:380247
n: 22 y:296877
n: 23 y:295944
n: 24 y:393028
n: 25 y:396226
n: 26 y:503947
n: 27 y:295944
n: 28 y:408831
n: 29 y:297410
n: 30 y:297571
n: 31 y:297009
n: 32 y:298164
n: 33 y:296247
n: 34 y:295944
n: 35 y:296688
n: 36 y:298019
n: 37 y:446420
n: 38 y:296757
n: 39 y:300672
n: 40 y:297820
n: 41 y:296726
n: 42 y:464563
n: 43 y:297132
n: 44 y:299200
n: 45 y:299218
n: 46 y:486119
n: 47 y:299288
n: 48 y:492852
n: 49 y:301054
n: 50 y:500010
n: 51 y:302702
n: 52 y:509514
n: 53 y:513044
n: 54 y:735044
n: 55 y:742565
n: 56 y:1198288
n: 57 y:2124530
n: 58 y:2157065
n: 59 y:2188002
n: 60 y:2222605
n: 61 y:2742437
n: 62 y:2781226
n: 63 y:2570251
n: 64 y:2860434
n: 65 y:2640806
n: 66 y:2941900
n: 67 y:2714345
n: 68 y:3021630
n: 69 y:3062854
n: 70 y:2820324
n: 71 y:2856964
n: 72 y:3182468
n: 73 y:3222512
n: 74 y:3262409
n: 75 y:3302960
n: 76 y:3343360
n: 77 y:3381396
n: 78 y:3421944
n: 79 y:3463492
n: 80 y:3501279
n: 81 y:3540978
n: 82 y:3581028
n: 83 y:3621288
n: 84 y:3660580
n: 85 y:3701580
n: 86 y:3742551
n: 87 y:3778856
n: 88 y:3821967
n: 89 y:3862207
n: 90 y:3903901
n: 91 y:3942269
n: 92 y:3982405
n: 93 y:4022748
n: 94 y:4062035
n: 95 y:4101398
n: 96 y:4143395
n: 97 y:4182780
n: 98 y:4222460
n: 99 y:4260776
n: 0 y:303273
n: 1 y:339788
n: 2 y:382334
n: 3 y:420801
n: 4 y:461949
n: 5 y:502981
n: 6 y:541944
n: 7 y:580836
n: 8 y:620034
n: 9 y:658923
n: 10 y:700888
n: 11 y:741252
n: 12 y:442780
n: 13 y:297302
n: 14 y:296757
n: 15 y:296898
n: 16 y:296617
n: 17 y:297258
n: 18 y:296350
n: 19 y:296108
n: 20 y:297414
n: 21 y:296722
n: 22 y:296332
n: 23 y:297400
n: 24 y:298321
n: 25 y:296932
n: 26 y:297444
n: 27 y:295944
n: 28 y:297710
n: 29 y:296980
n: 30 y:295944
n: 31 y:295944
n: 32 y:296712
n: 33 y:297414
n: 34 y:297476
n: 35 y:298116
n: 36 y:295944
n: 37 y:297852
n: 38 y:295944
n: 39 y:295944
n: 40 y:456236
n: 41 y:952319
n: 42 y:1135952
n: 43 y:295944
n: 44 y:647947
n: 45 y:476686
n: 46 y:664724
n: 47 y:486029
n: 48 y:1063950
n: 49 y:1668504
n: 50 y:1696628
n: 51 y:1724930
n: 52 y:1336333
n: 53 y:1779955
n: 54 y:1807955
n: 55 y:1175950
n: 56 y:2313066
n: 57 y:2349120
n: 58 y:1920828
n: 59 y:2183956
n: 60 y:1735953
n: 61 y:2491958
n: 62 y:2776544
n: 63 y:2563958
n: 64 y:2600704
n: 65 y:2636772
n: 66 y:2935960
n: 67 y:2708413
n: 68 y:3016961
n: 69 y:2782264
n: 70 y:2818663
n: 71 y:3137596
n: 72 y:3179407
n: 73 y:3216788
n: 74 y:3257054
n: 75 y:3295960
n: 76 y:3336700
n: 77 y:3375960
n: 78 y:3416612
n: 79 y:3457659
n: 80 y:3497452
n: 81 y:3537599
n: 82 y:3577268
n: 83 y:3616664
n: 84 y:3656240
n: 85 y:3695960
n: 86 y:3737040
n: 87 y:3776415
n: 88 y:3817015
n: 89 y:3856330
n: 90 y:3896700
n: 91 y:3936651
n: 92 y:3975960
n: 93 y:4015960
n: 94 y:4057728
n: 95 y:4095960
n: 96 y:4135960
n: 97 y:4177005
n: 98 y:4216401
n: 99 y:4255960
n: 0 y:303090
n: 1 y:343207
n: 2 y:382058
n: 3 y:422000
n: 4 y:463169
n: 5 y:503169
n: 6 y:541875
n: 7 y:581575
n: 8 y:621667
n: 9 y:660794
n: 10 y:701228
n: 11 y:698067
n: 12 y:734812
n: 13 y:300703
n: 14 y:354563
n: 15 y:300301
n: 16 y:300609
n: 17 y:299843
n: 18 y:299596
n: 19 y:299122
n: 20 y:300750
n: 21 y:299134
n: 22 y:299694
n: 23 y:301986
n: 24 y:299066
n: 25 y:299305
n: 26 y:300173
n: 27 y:300580
n: 28 y:300774
n: 29 y:297735
n: 30 y:299444
n: 31 y:300355
n: 32 y:299367
n: 33 y:298436
n: 34 y:297759
n: 35 y:298926
n: 36 y:301298
n: 37 y:299290
n: 38 y:299886
n: 39 y:298256
n: 40 y:298994
n: 41 y:299854
n: 42 y:299133
n: 43 y:299596
n: 44 y:300086
n: 45 y:300790
n: 46 y:299499
n: 47 y:300146
n: 48 y:298642
n: 49 y:299875
n: 50 y:499866
n: 51 y:302122
n: 52 y:301457
n: 53 y:726060
n: 54 y:1380889
n: 55 y:1621125
n: 56 y:972234
n: 57 y:1669504
n: 58 y:2158926
n: 59 y:2189500
n: 60 y:1981596
n: 61 y:2741047
n: 62 y:2530752
n: 63 y:2568061
n: 64 y:2860366
n: 65 y:2902683
n: 66 y:2413299
n: 67 y:2711514
n: 68 y:3020137
n: 69 y:3060779
n: 70 y:3102137
n: 71 y:3140295
n: 72 y:3180500
n: 73 y:2928128
n: 74 y:2965079
n: 75 y:3300054
n: 76 y:3342783
n: 77 y:3380688
n: 78 y:3422371
n: 79 y:3459906
n: 80 y:3502238
n: 81 y:3541903
n: 82 y:3581946
n: 83 y:3620914
n: 84 y:3662731
n: 85 y:3701584
n: 86 y:3741858
n: 87 y:3781074
n: 88 y:3822619
n: 89 y:3861918
n: 90 y:3900070
n: 91 y:3942786
n: 92 y:3981390
n: 93 y:4022870
n: 94 y:4059225
n: 95 y:4103278
n: 96 y:4141877
n: 97 y:4183108
n: 98 y:4220188
n: 99 y:4261345
n: 0 y:300650
n: 1 y:343242
n: 0 y:301046
n: 1 y:342904
n: 2 y:382428
n: 0 y:303888
n: 1 y:343856
n: 2 y:384040
